module ring_oscillator (reg vout);
output vout;
endmodule
