module adc1bit (reg in1, reg in2, reg out);
input in1;
input in2;
output out;
endmodule
